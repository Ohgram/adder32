program test;
    // typedef enum {IDLE,TEST,START} state;
    // enum bit[2:0]{S0='b001,S1='b010,S2='b100} st;
    // state c_st,n_st=IDLE;
    // $display( "st= %3b,n_st = %s",st,n_st.name);
    initial begin
    $display("hello,world");   
    end
    
endprogram